`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2022/03/10 18:53:45
// Design Name: 
// Module Name: exp_3
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module exp_3(
    output [3:0] q,
    input clk,
    input reset
    );

wire clk_1hz;
    
fre_divider_50M U0(.clk(clk), .reset(reset), .clk_new(clk_1hz));
exp_3_pre U1(.clk(clk_1hz), .reset(reset), .o(q));

endmodule
